// Custom defined datatypes

package types_pkg;

  typedef enum {
    READ,
    WRITE,
    EXECUTE
  } access_type_t;
 
 endpackage : types_pkg