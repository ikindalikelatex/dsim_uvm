package parameters_pkg;
  import types_pkg::*;

  // Define parameters for the adder
  parameter int ADDER_DATA_WIDTH = 8;
  parameter int COVERAGE_NUM_AUTO_BINS = 8;

endpackage : parameters_pkg