`include "uvm_macros.svh"

package sequences_pkg;
  // Import necessary UVM packages
  import uvm_pkg::*;
  import types_pkg::*;
  import parameters_pkg::*;
  import sequence_item_pkg::*;

  `include "base_sequence.sv"

endpackage : sequences_pkg