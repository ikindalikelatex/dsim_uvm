`include "uvm_macros.svh"

package env_pkg;
  import uvm_pkg::*;
  import types_pkg::*;
  import parameters_pkg::*;
  import agent_pkg::*;

  `include "environment.sv"
endpackage : env_pkg