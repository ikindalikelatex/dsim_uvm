`include "uvm_macros.svh"

package sequence_item_pkg;
  import uvm_pkg::*;
  import types_pkg::*;
  import parameters_pkg::*;

  `include "base_transaction.sv"
endpackage : sequence_item_pkg