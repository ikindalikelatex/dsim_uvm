package dpi_scoreboard_pkg;

  import "DPI-C" function longint unsigned dpi_get_sum(
    input longint unsigned a,
    input longint unsigned b
  );

endpackage : dpi_scoreboard_pkg