`include "uvm_macros.svh"

package test_pkg;
  import uvm_pkg::*;
  import types_pkg::*;
  import parameters_pkg::*;
  import sequence_item_pkg::*;
  import sequences_pkg::*;
  import env_pkg::*;

  `include "base_test.sv"
endpackage : test_pkg